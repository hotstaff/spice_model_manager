* JFET IV Curve Simulation
VDS 1 0 DC 0
VGS 2 0 DC 0
J1 1 2 0 2sk208

* JFET Model Parameters
.model 2SK208 NJF Vto=-2.638 Beta=1.059m Lambda=2.8m Rs=56.63 Rd=56.63 Betatce=-.5  Vtotc=-2.5m Cgd=10.38p M=.4373 Pb=.3905 Fc=.5 Cgs=6.043p Isr=112.8p Nr=2 Is=11.28p N=1 Xti=3 Alpha=10u Vk=100 Kf=1E-18

* DC Sweep for VDS with VGS as a parameter
.DC VDS 0 20 0.1 VGS -0.4 0 0.1

* Output the data to file
.control
    run
    set wr_vecnames
    wrdata /home/hotstaff/spice_model_manager/simulation/data/jfet_iv_curve_data.dat V(1) I(VDS) V(2)  ; V(2)はVGSを出力
.endc

.print DC V(1) I(VDS) V(2)

.end